package orion_soc_types;
    // parameter SOC_IMEM_SIZE = 32*1024;   // 32KB
    // parameter SOC_DMEM_SIZE = 32*1024;   // 32KB  

    parameter SOC_MEM_ADDR = 32'h0001_0000;
    parameter SOC_MEM_SIZE = 64*1024;       // 64KB
endpackage
