package orion_soc_types;
    parameter SOC_IMEM_SIZE = 32*1024;     // 32KB
    parameter SOC_DMEM_SIZE = 32*1024;     // 32KB  
endpackage
